--BCD Counter Entity
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY BCD_CNT IS
	PORT ( CLK : IN  STD_LOGIC;
		RESET : IN  STD_LOGIC;
		DOUT12 : OUT  STD_LOGIC_VECTOR (11 DOWNTO 0)
	);
END ENTITY BCD_CNT;

ARCHITECTURE ART1 OF BCD_CNT IS
	SIGNAL BCD_CNT_REG : STD_LOGIC_VECTOR(11 DOWNTO 0);
BEGIN
	PROCESS(CLK)
	BEGIN
		IF(CLK'EVENT AND CLK='1') THEN
			DOUT12 <= BCD_CNT_REG;
		END IF;	
	END PROCESS;
	PROCESS(CLK,RESET)
	BEGIN
		IF RESET = '0' THEN
			BCD_CNT_REG(3 DOWNTO 0) <= (OTHERS=> '0');
		ELSIF(CLK'EVENT AND CLK='1') THEN
			--低4位遇9变0
			IF (BCD_CNT_REG(3 DOWNTO 0) = "1001") THEN
				BCD_CNT_REG(3 DOWNTO 0) <= (OTHERS=> '0');
			ELSE
				BCD_CNT_REG(3 DOWNTO 0) <= BCD_CNT_REG(3 DOWNTO 0) + 1;
			END IF;
		END IF;
	END PROCESS;
	
	PROCESS(CLK,RESET)
	BEGIN
		IF RESET = '0' THEN
		BCD_CNT_REG(7 DOWNTO 4) <= (OTHERS=> '0');
	ELSIF(CLK'EVENT AND CLK='1') THEN
		--中间4位先判断是否有低4位的进位，有才会计数
		IF (BCD_CNT_REG(3 DOWNTO 0) = "1001") THEN
			IF (BCD_CNT_REG(7 DOWNTO 4) = "1001") THEN
				BCD_CNT_REG(7 DOWNTO 4) <= (OTHERS=> '0');
			ELSE
				BCD_CNT_REG(7 DOWNTO 4) <= BCD_CNT_REG(7 DOWNTO 4) + 1;
			END IF;
		ELSE
			BCD_CNT_REG(7 DOWNTO 4) <= BCD_CNT_REG(7 DOWNTO 4);
		END IF;
	END IF;
	END PROCESS;
	
	PROCESS(CLK,RESET)
	BEGIN
		IF RESET = '0' THEN
			BCD_CNT_REG(11 DOWNTO 8) <= (OTHERS=> '0');
		ELSIF(CLK'EVENT AND CLK='1') THEN
		--高4位先判断是否有来自中间4位的进位
			IF (BCD_CNT_REG(7 DOWNTO 4) = "1001") THEN
				IF (BCD_CNT_REG(11 DOWNTO 8) = "1001") THEN
					BCD_CNT_REG(11 DOWNTO 8) <= (OTHERS=> '0');
				ELSE
					BCD_CNT_REG(11 DOWNTO 8) <= BCD_CNT_REG(11 DOWNTO 8) + 1;
				END IF;
			ELSE
				BCD_CNT_REG(11 DOWNTO 8) <= BCD_CNT_REG(11 DOWNTO 8);
			END IF;
		END IF;
	END PROCESS;  
END ARCHITECTURE ART1;