--4选1数据选择器
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
ENTITY MUXB41 IS
	PORT(DATA0,DATA1,DATA2,DATA3:IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		A,B:IN STD_LOGIC;
		Y:OUT STD_LOGIC_VECTOR(3 DOWNTO 0));
END ENTITY;		
ARCHITECTURE ART OF MUXB41 IS
	SIGNAL SEL:STD_LOGIC_VECTOR(1 DOWNTO 0);
	BEGIN
	SEL<=B&A;
	PROCESS(SEL)
		BEGIN
		CASE SEL IS
			WHEN "00"=>Y<=DATA0;
			WHEN "01"=>Y<=DATA1;
			WHEN "10"=>Y<=DATA2;
			WHEN "11"=>Y<=DATA3;
			WHEN OTHERS=>Y<=NULL;
		END CASE;
	END PROCESS;
END ARCHITECTURE ART;