--Led Display
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY LED_DISP IS
PORT(	CLK_DISP		:IN 	STD_LOGIC;
		DATA_IN_1	:IN 	STD_LOGIC_VECTOR(3 DOWNTO 0);
		DATA_IN_2	:IN 	STD_LOGIC_VECTOR(3 DOWNTO 0);
		DATA_IN_3	:IN 	STD_LOGIC_VECTOR(3 DOWNTO 0);
		DATA2LED		:OUT 	STD_LOGIC_VECTOR(6 DOWNTO 0);
		SEL2LED		:OUT 	STD_LOGIC_VECTOR(2 DOWNTO 0));

END ENTITY LED_DISP;

ARCHITECTURE ART1 OF LED_DISP IS
SIGNAL DOUT_OCT: STD_LOGIC_VECTOR (3 DOWNTO 0);
BEGIN
	PROCESS (CLK_DISP)
		VARIABLE VAR: STD_LOGIC_VECTOR (1 DOWNTO 0):="00";
		
		BEGIN	
			IF(CLK_DISP 'EVENT AND CLK_DISP='1') THEN
				IF(VAR="11")THEN 
					VAR:="00";
				END IF;	
				IF(VAR="00")THEN
					SEL2LED <="001";
					DOUT_OCT <= DATA_IN_1;
				ELSIF(VAR="01")THEN
					SEL2LED <="010";
					DOUT_OCT <= DATA_IN_2;
				ELSE
					SEL2LED <="100";
					DOUT_OCT <= DATA_IN_3;
				END IF;
				VAR:=VAR+1;							
			END IF;							
	END PROCESS;
	PROCESS(DOUT_OCT)
	BEGIN
		CASE DOUT_OCT IS
			WHEN"0000"=> DATA2LED <="1111110";
			WHEN"0001"=> DATA2LED <="0110000";
			WHEN"0010"=> DATA2LED <="1101101";
			WHEN"0011"=> DATA2LED <="1111001";
			WHEN"0100"=> DATA2LED <="0110011";
			WHEN"0101"=> DATA2LED <="1011011";
			WHEN"0110"=> DATA2LED <="1011111";
			WHEN"0111"=> DATA2LED <="1110000";
			WHEN"1000"=> DATA2LED <="1111111";
			WHEN"1001"=> DATA2LED <="1111011";
			WHEN OTHERS => DATA2LED <="0000000";
		END CASE;	
	END PROCESS;		
END ARCHITECTURE ART1;

