--Select Signal
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY SEL_SIGNAL IS
PORT(
		TEST_CLK		:IN STD_LOGIC;
		MEASURE_CLK	:IN STD_LOGIC;
		CHOOSE		:IN STD_LOGIC;
		CLK			:OUT STD_LOGIC);

END ENTITY SEL_SIGNAL;

ARCHITECTURE ART1 OF SEL_SIGNAL IS
	BEGIN 
	PROCESS(TEST_CLK,MEASURE_CLK,CHOOSE)
		BEGIN
		IF (CHOOSE='0') THEN
			CLK<=TEST_CLK;
		ELSE
			CLK<=MEASURE_CLK;
		END IF;
	END PROCESS;

END ART1;

