LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
--自定义程序包
PACKAGE MYTYPE IS
SUBTYPE PIXEL IS INTEGER RANGE 0 TO 255;
TYPE MATRIX IS ARRAY(0 TO 255, 0 TO 255) OF INTEGER;
END PACKAGE MYTYPE;
PACKAGE BODY MYTYPE IS
END MYTYPE;