LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
ENTITY CHKSEQ IS
	PORT(DIN:IN STD_LOGIC;
		  CLK,RESET:IN STD_LOGIC;
		  DOUT:OUT STD_LOGIC);
END ENTITY CHKSEQ;
ARCHITECTURE ART OF CHKSEQ IS
	TYPE STATETYPE IS(S1,S2,S3,S4,S5,S6,S7,S8);
	SIGNAL PRESENT_STATE,NEXT_STATE:STATETYPE;
BEGIN
	COMB_PROCESS:PROCESS(DIN,PRESENT_STATE)
	BEGIN
		CASE PRESENT_STATE IS
			WHEN S1=>DOUT<='0';
				IF DIN='0' THEN
					NEXT_STATE<=S1;
				ELSE
					NEXT_STATE<=S2;
				END IF;
			WHEN S2=>DOUT<='0';
				IF DIN='0' THEN
					NEXT_STATE<=S2;
				ELSE
					NEXT_STATE<=S3;
				END IF;
			WHEN S3=>DOUT<='0';
				IF DIN='0' THEN
					NEXT_STATE<=S1;
				ELSE
					NEXT_STATE<=S4;
				END IF;
			WHEN S4=>DOUT<='0';
				IF DIN='0' THEN
					NEXT_STATE<=S5;
				ELSE
					NEXT_STATE<=S4;
				END IF;
			WHEN S5=>DOUT<='0';
				IF DIN='0' THEN
					NEXT_STATE<=S6;
				ELSE
					NEXT_STATE<=S2;
				END IF;
			WHEN S6=>DOUT<='0';
				IF DIN='0' THEN
					NEXT_STATE<=S1;
				ELSE
					NEXT_STATE<=S7;
				END IF;
			WHEN S7=>DOUT<='0';
				IF DIN='0' THEN
					NEXT_STATE<=S8;
				ELSE
					NEXT_STATE<=S3;
				END IF;
			WHEN S8=>DOUT<='1';
				IF DIN='0' THEN
					NEXT_STATE<=S1;
				ELSE
					NEXT_STATE<=S2;
				END IF;
		END CASE;		
	END PROCESS;
	
	CLK_PROCESS:PROCESS(CLK,RESET)
	BEGIN
		IF(RESET='1') THEN
			PRESENT_STATE<=S1;
		ELSIF(CLK'EVENT AND CLK='1') THEN
			PRESENT_STATE<=NEXT_STATE;
		END IF;
	END PROCESS;
END ARCHITECTURE ART;	