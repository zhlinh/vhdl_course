--LED Decoder Entity
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY LED_DEC IS
	PORT ( NUM : IN  STD_LOGIC_VECTOR (3 DOWNTO 0);
			DOUT : OUT  STD_LOGIC_VECTOR (6 DOWNTO 0)
	);
END ENTITY LED_DEC;

ARCHITECTURE ART1 OF LED_DEC IS
BEGIN
	PROCESS(NUM)
	BEGIN
		CASE(NUM) IS
			WHEN "0000" =>
				DOUT <= "1111110";
			WHEN "0001" =>
				DOUT <= "0110000";
			WHEN "0010" =>
				DOUT <= "1101101";
			WHEN "0011" =>
				DOUT <= "1111001";
			WHEN "0100" =>
				DOUT <= "0110011";
			WHEN "0101" =>
				DOUT <= "1011011";
			WHEN "0110" =>
				DOUT <= "1011111";
			WHEN "0111" =>
				DOUT <= "1110000";
			WHEN "1000" =>
				DOUT <= "1111111";
			WHEN "1001" =>
				DOUT <= "1111011";
			WHEN OTHERS =>
				DOUT <= (OTHERS=> '0');
		END CASE;
	END PROCESS;
END ARCHITECTURE ART1;