--Top Entity
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY FREQ_CNT IS
PORT(
		RST:              IN STD_LOGIC;
		CLK_IN_1HZ:       IN STD_LOGIC;
		CLK_DISP:         IN STD_LOGIC;
		TEST_CLK:         IN STD_LOGIC;
		MEASURE_CLK:      IN STD_LOGIC;
		CHOOSE:           IN STD_LOGIC;
		DATA_RANGE:       IN STD_LOGIC;

		BEEP:             OUT STD_LOGIC;
		RANGE_DISP:       OUT STD_LOGIC;
		DATA2LED:         OUT 	STD_LOGIC_VECTOR(6 DOWNTO 0);
		SEL2LED:          OUT 	STD_LOGIC_VECTOR(2 DOWNTO 0));

END ENTITY FREQ_CNT;



ARCHITECTURE ART OF FREQ_CNT IS

	COMPONENT DIV_FREQ IS
	PORT(	CLK_IN_1HZ:   IN STD_LOGIC;
			RST:          IN STD_LOGIC;
			CLK_OUT_05HZ: OUT STD_LOGIC);
	END COMPONENT;

	COMPONENT SEL_SIGNAL IS
	PORT(	TEST_CLK:     IN STD_LOGIC;
			MEASURE_CLK:  IN STD_LOGIC;
			CHOOSE:       IN STD_LOGIC;
			CLK:          OUT STD_LOGIC);
	END COMPONENT;

	COMPONENT COUNT IS
	PORT(	CLK:          IN 	STD_LOGIC;
			CLK_OUT_05HZ: IN 	STD_LOGIC;
			RST:          IN 	STD_LOGIC;
			D1:           OUT 	STD_LOGIC_VECTOR(3 DOWNTO 0);
			D2:           OUT 	STD_LOGIC_VECTOR(3 DOWNTO 0);
			D3:           OUT 	STD_LOGIC_VECTOR(3 DOWNTO 0);
			D4:           OUT 	STD_LOGIC_VECTOR(3 DOWNTO 0);
			CARRY:        OUT 	STD_LOGIC;
			READ_EN:      OUT	STD_LOGIC);
	END COMPONENT;

	COMPONENT ALERT IS
	PORT(	DATA_RANGE:   IN STD_LOGIC;
			CARRY_LABEL:  IN STD_LOGIC;
			D1_IN:        IN STD_LOGIC_VECTOR(3 DOWNTO 0);
			D2_IN:        IN STD_LOGIC_VECTOR(3 DOWNTO 0);
			D3_IN:        IN STD_LOGIC_VECTOR(3 DOWNTO 0);
			D4_IN:        IN STD_LOGIC_VECTOR(3 DOWNTO 0);

			D1_OUT:       OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
			D2_OUT:       OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
			D3_OUT:       OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
			BEEP:         OUT STD_LOGIC;
			RANGE_DISP:   OUT STD_LOGIC);
	END COMPONENT;

	COMPONENT D_LATCH IS
	PORT(	LATCH_EN:     IN STD_LOGIC;
			D1_IN:        IN STD_LOGIC_VECTOR(3 DOWNTO 0);
			D2_IN:        IN STD_LOGIC_VECTOR(3 DOWNTO 0);
			D3_IN:        IN STD_LOGIC_VECTOR(3 DOWNTO 0);
			D1_OUT:       OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
			D2_OUT:       OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
			D3_OUT:       OUT STD_LOGIC_VECTOR(3 DOWNTO 0));
	END COMPONENT;

	COMPONENT LED_DISP IS
	PORT(	CLK_DISP:     IN STD_LOGIC;
			DATA_IN_1:    IN STD_LOGIC_VECTOR(3 DOWNTO 0);
			DATA_IN_2:    IN STD_LOGIC_VECTOR(3 DOWNTO 0);
			DATA_IN_3:    IN STD_LOGIC_VECTOR(3 DOWNTO 0);
			DATA2LED:     OUT STD_LOGIC_VECTOR(6 DOWNTO 0);
			SEL2LED:      OUT STD_LOGIC_VECTOR(2 DOWNTO 0));
	END COMPONENT;


	SIGNAL WIRE1:         STD_LOGIC;
	SIGNAL WIRE2:         STD_LOGIC;
	SIGNAL WIRE3:         STD_LOGIC;
	SIGNAL WIRE4:         STD_LOGIC;
	SIGNAL WIRE_C_D1:     STD_LOGIC_VECTOR(3 DOWNTO 0);
	SIGNAL WIRE_C_D2:     STD_LOGIC_VECTOR(3 DOWNTO 0);
	SIGNAL WIRE_C_D3:     STD_LOGIC_VECTOR(3 DOWNTO 0);
	SIGNAL WIRE_C_D4:     STD_LOGIC_VECTOR(3 DOWNTO 0);

	SIGNAL WIRE_A_D1:     STD_LOGIC_VECTOR(3 DOWNTO 0);
	SIGNAL WIRE_A_D2:     STD_LOGIC_VECTOR(3 DOWNTO 0);
	SIGNAL WIRE_A_D3:     STD_LOGIC_VECTOR(3 DOWNTO 0);

	SIGNAL WIRE_L_D1:     STD_LOGIC_VECTOR(3 DOWNTO 0);
	SIGNAL WIRE_L_D2:     STD_LOGIC_VECTOR(3 DOWNTO 0);
	SIGNAL WIRE_L_D3:     STD_LOGIC_VECTOR(3 DOWNTO 0);

	BEGIN
	INST_DIV_FREQ:       DIV_FREQ
		PORT MAP(CLK_IN_1HZ      => CLK_IN_1HZ,
					RST          => RST,
					CLK_OUT_05HZ => WIRE1);


	INST_SEL_SIGNAL:      SEL_SIGNAL
		PORT MAP(TEST_CLK        => TEST_CLK,
					MEASURE_CLK  => MEASURE_CLK,
					CHOOSE       => CHOOSE,
					CLK          => WIRE2);

	INST_COUNT:         COUNT
		PORT MAP(CLK             => WIRE2,
					CLK_OUT_05HZ => WIRE1,
					RST          => RST,
					D1           => WIRE_C_D1,
					D2           => WIRE_C_D2,
					D3           => WIRE_C_D3,
					D4           => WIRE_C_D4,
					CARRY        => WIRE3,
					READ_EN      => WIRE4);

	INST_ALERT:           ALERT
		PORT MAP(DATA_RANGE      => DATA_RANGE,
					CARRY_LABEL  => WIRE3,
					D1_IN        => WIRE_C_D1,
					D2_IN        => WIRE_C_D2,
					D3_IN        => WIRE_C_D3,
					D4_IN        => WIRE_C_D4,
					D1_OUT       => WIRE_A_D1,
					D2_OUT       => WIRE_A_D2,
					D3_OUT       => WIRE_A_D3,
					BEEP         => BEEP,
					RANGE_DISP   => RANGE_DISP);

	INST_D_LATCH:           D_LATCH
		PORT MAP(LATCH_EN        => WIRE4,
					D1_IN        => WIRE_A_D1,
					D2_IN        => WIRE_A_D2,
					D3_IN        => WIRE_A_D3,
					D1_OUT       => WIRE_L_D1,
					D2_OUT       => WIRE_L_D2,
					D3_OUT       => WIRE_L_D3);

	INST_LED_DISP:        LED_DISP
		PORT MAP(CLK_DISP        => CLK_DISP,
					DATA_IN_1    => WIRE_L_D1,
					DATA_IN_2    => WIRE_L_D2,
					DATA_IN_3    => WIRE_L_D3,
					DATA2LED     => DATA2LED,
					SEL2LED      => SEL2LED);

END ARCHITECTURE ART;

