--4选1信号选择器
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
ENTITY MUX41 IS
	PORT(X:IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		A,B:IN STD_LOGIC;
		Y:OUT STD_LOGIC);
END ENTITY MUX41;
ARCHITECTURE ART OF MUX41 IS
	SIGNAL SEL:STD_LOGIC_VECTOR(1 DOWNTO 0);
	BEGIN
	SEL<=B&A;
	PROCESS(X,SEL) IS
		BEGIN
		IF(SEL="00") THEN Y<=X(0);
		ELSIF(SEL="01") THEN Y<=X(1);
		ELSIF(SEL="11") THEN Y<=X(2);
		ELSE Y<=X(3);
		END IF;
	END PROCESS;
END ARCHITECTURE ART;