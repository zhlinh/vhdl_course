--Frequency Divider
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY DIV_FREQ IS
	PORT(	CLK_IN_1HZ	:IN STD_LOGIC;
			RST			:IN STD_LOGIC;
			CLK_OUT_05HZ:OUT STD_LOGIC);
END ENTITY DIV_FREQ;


ARCHITECTURE ART1 OF DIV_FREQ IS

	BEGIN
	PROCESS (CLK_IN_1HZ,RST)
	VARIABLE  CLK_OUT_TEMP:STD_LOGIC_VECTOR (1 DOWNTO 0):="00";
		BEGIN
		IF(RST='1')THEN
			CLK_OUT_TEMP:="00";
			ELSE IF(CLK_IN_1HZ 'EVENT AND CLK_IN_1HZ='1')THEN
				CLK_OUT_TEMP := CLK_OUT_TEMP + "01";
			END IF;
		END IF;
		CLK_OUT_05HZ <= CLK_OUT_TEMP(0);
	END PROCESS;

END ARCHITECTURE ART1;

