LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
ENTITY TB_CHKSEQ IS
END ENTITY TB_CHKSEQ;
ARCHITECTURE DIRECT_WAY OF TB_CHKSEQ IS
	COMPONENT CHKSEQ
		PORT(CLK,RESET,DIN:IN STD_LOGIC;
			 DOUT:OUT STD_LOGIC);
	END COMPONENT;
SIGNAL CLK,RESET,DIN:STD_LOGIC:='0';
SIGNAL 	DOUT:STD_LOGIC;
SIGNAL	GIVEN_SEQ:STD_LOGIC_VECTOR(48 DOWNTO 0)
				 :="0111110010010110111011011101110111111100101110010";
CONSTANT CLK_PERIOD:TIME:=10 NS;
BEGIN
-- DUT = DEVICE UNDER TEST
	DUT:CHKSEQ PORT MAP(
			CLK=>CLK,
			RESET=>RESET,
			DIN=>DIN,
			DOUT=>DOUT);
--CLOCK PROCESS
	CLK_PROCESS:PROCESS
	BEGIN
		CLK<='0';
		WAIT FOR CLK_PERIOD/2;
		CLK<='1';
		WAIT FOR CLK_PERIOD/2;
	END PROCESS;
--GIVEN SEQUENCE PROCESS
	GIVEN_SEQ_PROCESS:PROCESS(CLK)
	BEGIN
		
		IF(CLK'EVENT AND CLK='1') THEN
			GIVEN_SEQ<=GIVEN_SEQ(47 DOWNTO 0) & '0';
			DIN<=GIVEN_SEQ(48);
		END IF;
	END PROCESS;
--SET UP THE RESET SIGNAL
	STIMULIS_PROCESS:PROCESS 
	BEGIN
		RESET<='1';
		WAIT FOR CLK_PERIOD;
		RESET<='0';
		WAIT FOR CLK_PERIOD*8;
		RESET<='1';
		WAIT FOR CLK_PERIOD/2;
		RESET<='0';
		WAIT;
	END	PROCESS;
END ARCHITECTURE DIRECT_WAY;	
		
