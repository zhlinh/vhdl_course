--Top-Level Entity
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY LED_CNT IS 
	PORT ( 
		CLK : IN  STD_LOGIC; ---THE CLK OF CNT
	   CLKDSP : IN  STD_LOGIC; ---THE CLK OF SACN
	   RESET : IN  STD_LOGIC;
	   DOUT : OUT  STD_LOGIC_VECTOR (6 DOWNTO 0);
	   SEL : OUT  STD_LOGIC_VECTOR (1 DOWNTO 0)
	);
END ENTITY LED_CNT;

ARCHITECTURE ART OF LED_CNT IS

	COMPONENT BCD_CNT
	PORT(
		CLK : IN STD_LOGIC;
		RESET : IN STD_LOGIC;
		DOUT12 : OUT STD_LOGIC_VECTOR(11 DOWNTO 0)
	);
	END COMPONENT;

	COMPONENT SCANNER
	PORT(
		CLK_SCAN : IN STD_LOGIC;
		RESET : IN STD_LOGIC;
		DIN12 : IN STD_LOGIC_VECTOR(11 DOWNTO 0);          
		NUM : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		SEL : OUT STD_LOGIC_VECTOR(1 DOWNTO 0)
	);
	END COMPONENT;
	
	COMPONENT LED_DEC
	PORT(
		NUM : IN STD_LOGIC_VECTOR(3 DOWNTO 0);          
		DOUT : OUT STD_LOGIC_VECTOR(6 DOWNTO 0)
	);
	END COMPONENT;
	
	SIGNAL BCD_CNT_MID1 : STD_LOGIC_VECTOR(11 DOWNTO 0);
	SIGNAL SCAN_MID2 : STD_LOGIC_VECTOR(3 DOWNTO 0);
	
BEGIN
	INST_BCD_CNT : BCD_CNT PORT MAP(
		CLK => CLK,
		RESET => RESET,
		DOUT12 => BCD_CNT_MID1
	);
	INST_SCANNER : SCANNER PORT MAP(
		CLK_SCAN => CLKDSP,
		RESET => RESET,
		DIN12 => BCD_CNT_MID1,
		NUM => SCAN_MID2,
		SEL => SEL
	);
  	INST_LED_DEC: LED_DEC PORT MAP(
		NUM => SCAN_MID2,
		DOUT => DOUT
	);
END ARCHITECTURE ART;