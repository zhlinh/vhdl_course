--比较两个二进制数是否相等
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
ENTITY COMPARE IS
	PORT(A,B:IN STD_LOGIC_VECTOR(7 DOWNTO 0);
			EQ:OUT STD_LOGIC);
END ENTITY COMPARE;
ARCHITECTURE ART OF COMPARE IS
	BEGIN
	EQ<='1' WHEN A=B ELSE '0';
END ARCHITECTURE ART;	