--MYTYPE package
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
--自定义程序包
PACKAGE MYTYPE IS
    SUBTYPE COLOR IS INTEGER RANGE 0 TO 255;
    FUNCTION CONV_TO_CHAR   (SLV8 :STD_LOGIC_VECTOR (7 DOWNTO 0)) RETURN CHARACTER;
    FUNCTION CONV_TO_VECTOR   (CHAR :CHARACTER)  RETURN STD_LOGIC_VECTOR;
END PACKAGE MYTYPE;
PACKAGE BODY MYTYPE IS
    FUNCTION CONV_TO_CHAR (SLV8 :STD_LOGIC_VECTOR (7 DOWNTO 0)) RETURN CHARACTER IS
    CONSTANT XMAP :INTEGER :=0;
    VARIABLE TEMP :INTEGER :=0;
    BEGIN
        FOR I IN SLV8'RANGE LOOP
            TEMP:=TEMP*2;
            CASE SLV8(I) IS
                WHEN '0'   => NULL;
                WHEN '1'   => TEMP :=TEMP+1;
                WHEN OTHERS     => TEMP :=TEMP+XMAP;
            END CASE;
        END LOOP;
        RETURN CHARACTER'VAL(TEMP);
    END CONV_TO_CHAR;

    FUNCTION CONV_TO_VECTOR (CHAR :CHARACTER) RETURN STD_LOGIC_VECTOR IS
        VARIABLE SLV8 :STD_LOGIC_VECTOR (7 DOWNTO 0);
        VARIABLE TEMP :INTEGER :=CHARACTER'POS(CHAR);
    BEGIN
        FOR I IN SLV8'REVERSE_RANGE LOOP
            CASE TEMP MOD 2 IS
                WHEN 0 => SLV8(I):='0';
                WHEN 1 => SLV8(I):='1';
                WHEN OTHERS => NULL;
            END CASE;
            TEMP:=TEMP/2;
        END LOOP;
        RETURN SLV8;
    END CONV_TO_VECTOR;
END MYTYPE;
