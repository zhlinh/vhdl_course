LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
ENTITY TRISTATE IS
	PORT(EN,DIN:IN STD_LOGIC;
		DOUT:OUT STD_LOGIC);
END ENTITY TRISTATE;
ARCHITECTURE ART OF TRISTATE IS
	BEGIN
	PROCESS(EN,DIN) IS
		BEGIN
		IF EN='1' THEN
			DOUT<=DIN;
		ELSE
			DOUT<='Z';
		END IF;
	END PROCESS;
END ARCHITECTURE ART;