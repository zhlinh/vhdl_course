LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
ENTITY CHK_3BIT IS
	PORT(DIN:IN STD_LOGIC;
		CLK,RESET:IN STD_LOGIC;
		DOUT:OUT STD_LOGIC);
END ENTITY CHK_3BIT;  
ARCHITECTURE ART1 OF CHK_3BIT IS
	TYPE STATETYPE IS(S1,S2,S3,S4);
	SIGNAL PRESENT_STATE,NEXT_STATE:STATETYPE;
BEGIN
	COMB:PROCESS(PRESENT_STATE,DIN)
	BEGIN
		CASE PRESENT_STATE IS
			WHEN S1=>DOUT<='0';
				IF DIN='0'THEN
					NEXT_STATE<=S1;
				ELSE
					NEXT_STATE<=S2;
				END IF;
			WHEN S2=>DOUT<='0';
				IF DIN='0'THEN
					NEXT_STATE<=S1;
				ELSE
					NEXT_STATE<=S3;
				END IF;
			WHEN S3=>DOUT<='0';
				IF DIN='0'THEN
					NEXT_STATE<=S4;
				ELSE
					NEXT_STATE<=S3;
				END IF;
			WHEN S4=>DOUT<='1';
				IF DIN='0'THEN
					NEXT_STATE<=S1;
				ELSE
					NEXT_STATE<=S2;
				END IF;
		END CASE;
	END PROCESS;
	CLOCK:PROCESS(CLK,RESET)
	BEGIN
		IF(RESET='1')THEN
			PRESENT_STATE<=S1;
		ELSIF(CLK'EVENT AND CLK='1')THEN
			PRESENT_STATE<=NEXT_STATE;
		END IF;
	END PROCESS;
END ARCHITECTURE ART1;
