--Latch
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY D_LATCH IS
PORT(	LATCH_EN: IN STD_LOGIC;
		D1_IN:    IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		D2_IN:    IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		D3_IN:    IN STD_LOGIC_VECTOR(3 DOWNTO 0);

		D1_OUT:   OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		D2_OUT:   OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		D3_OUT:   OUT STD_LOGIC_VECTOR(3 DOWNTO 0));
END ENTITY D_LATCH;

ARCHITECTURE ART1 OF D_LATCH IS

BEGIN
	PROCESS(LATCH_EN)
	BEGIN
	 IF (LATCH_EN='1') THEN
		D1_OUT <= D1_IN;
		D2_OUT <= D2_IN;
		D3_OUT <= D3_IN;
	ELSE
		D1_OUT <= "0000";
		D2_OUT <= "0000";
		D3_OUT <= "0000";
	END IF;

	END PROCESS;
END ARCHITECTURE ART1;

