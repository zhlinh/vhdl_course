LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
ENTITY CHK_3BIT IS
	PORT(DIN:IN STD_LOGIC;
		CLK,RESET:IN STD_LOGIC;
		BIT3:IN STD_LOGIC_VECTOR(2 DOWNTO 0);
		DOUT:OUT STD_LOGIC);
END ENTITY CHK_3BIT;  
ARCHITECTURE ART1 OF CHK_3BIT IS
	TYPE STATETYPE IS(S1,S2,S3,S4,S5,S6,S7,S8,S9,S10,S11,S12,S13,S14,S15);
	SIGNAL PRESENT_STATE,NEXT_STATE:STATETYPE;
	SIGNAL CHOSEN_SEQ:STD_LOGIC_VECTOR(7 DOWNTO 0):="00000000";
BEGIN
	CHOOSE:PROCESS(BIT3)
	BEGIN
	--使用case语句时一定要列举完所有情况(善于应用others)，否则编译通过但仿真通不过
		CASE BIT3 IS
			WHEN "000"=>CHOSEN_SEQ<="00000001";
			WHEN "001"=>CHOSEN_SEQ<="00000010";
			WHEN "010"=>CHOSEN_SEQ<="00000100";
			WHEN "011"=>CHOSEN_SEQ<="00001000";
			WHEN "100"=>CHOSEN_SEQ<="00010000";
			WHEN "101"=>CHOSEN_SEQ<="00100000";
			WHEN "110"=>CHOSEN_SEQ<="01000000";
			WHEN "111"=>CHOSEN_SEQ<="10000000";
			WHEN OTHERS =>CHOSEN_SEQ<="00000000";
		END CASE;
	END PROCESS;	
	COMB:PROCESS(PRESENT_STATE,DIN)
	BEGIN
		CASE PRESENT_STATE IS
			WHEN S1=>DOUT<='0';
				IF DIN='0'THEN
					NEXT_STATE<=S2;
				ELSE
					NEXT_STATE<=S3;
				END IF;
			WHEN S2=>DOUT<='0';
				IF DIN='0'THEN
					NEXT_STATE<=S4;
				ELSE
					NEXT_STATE<=S5;
				END IF;
			WHEN S3=>DOUT<='0';
				IF DIN='0'THEN
					NEXT_STATE<=S6;
				ELSE
					NEXT_STATE<=S7;
				END IF;
			WHEN S4=>DOUT<='0';
				IF DIN='0'THEN
					NEXT_STATE<=S8;
				ELSE
					NEXT_STATE<=S9;
				END IF;
			WHEN S5=>DOUT<='0';
				IF DIN='0'THEN
					NEXT_STATE<=S10;
				ELSE
					NEXT_STATE<=S11;
				END IF;
			WHEN S6=>DOUT<='0';
				IF DIN='0'THEN
					NEXT_STATE<=S12;
				ELSE
					NEXT_STATE<=S13;
				END IF;
			WHEN S7=>DOUT<='0';
				IF DIN='0'THEN
					NEXT_STATE<=S14;
				ELSE
					NEXT_STATE<=S15;
				END IF;
			WHEN S8=>DOUT<=CHOSEN_SEQ(0);
				IF DIN='0'THEN
					NEXT_STATE<=S8;
				ELSE
					NEXT_STATE<=S9;
				END IF;
			WHEN S9=>DOUT<=CHOSEN_SEQ(1);
				IF DIN='0'THEN
					NEXT_STATE<=S10;
				ELSE
					NEXT_STATE<=S11;
				END IF;
			WHEN S10=>DOUT<=CHOSEN_SEQ(2);
				IF DIN='0'THEN
					NEXT_STATE<=S12;
				ELSE
					NEXT_STATE<=S13;
				END IF;
			WHEN S11=>DOUT<=CHOSEN_SEQ(3);
				IF DIN='0'THEN
					NEXT_STATE<=S14;
				ELSE
					NEXT_STATE<=S15;
				END IF;
			WHEN S12=>DOUT<=CHOSEN_SEQ(4);
				IF DIN='0'THEN
					NEXT_STATE<=S8;
				ELSE
					NEXT_STATE<=S9;
				END IF;
			WHEN S13=>DOUT<=CHOSEN_SEQ(5);
				IF DIN='0'THEN
					NEXT_STATE<=S10;
				ELSE
					NEXT_STATE<=S11;
				END IF;
			WHEN S14=>DOUT<=CHOSEN_SEQ(6);
				IF DIN='0'THEN
					NEXT_STATE<=S12;
				ELSE
					NEXT_STATE<=S13;
				END IF;
			WHEN S15=>DOUT<=CHOSEN_SEQ(7);
				IF DIN='0'THEN
					NEXT_STATE<=S14;
				ELSE
					NEXT_STATE<=S15;
				END IF;
		END CASE;
	END PROCESS;
	CLOCK:PROCESS(CLK,RESET)
	BEGIN
		IF(RESET='1')THEN
			PRESENT_STATE<=S1;
		ELSIF(CLK'EVENT AND CLK='1')THEN
			PRESENT_STATE<=NEXT_STATE;
		END IF;
	END PROCESS;
END ARCHITECTURE ART1;
